library verilog;
use verilog.vl_types.all;
entity Cache_sv_unit is
end Cache_sv_unit;
