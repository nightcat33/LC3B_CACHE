library verilog;
use verilog.vl_types.all;
entity Array_sv_unit is
end Array_sv_unit;
