library verilog;
use verilog.vl_types.all;
entity unadj_sv_unit is
end unadj_sv_unit;
