library verilog;
use verilog.vl_types.all;
entity nzp_sv_unit is
end nzp_sv_unit;
