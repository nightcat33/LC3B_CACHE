library verilog;
use verilog.vl_types.all;
entity sign_extend_sv_unit is
end sign_extend_sv_unit;
