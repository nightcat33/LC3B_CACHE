library verilog;
use verilog.vl_types.all;
entity CPU_sv_unit is
end CPU_sv_unit;
