library verilog;
use verilog.vl_types.all;
entity mp2 is
end mp2;
