library verilog;
use verilog.vl_types.all;
entity unsign_extend_sv_unit is
end unsign_extend_sv_unit;
