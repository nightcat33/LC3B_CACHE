library verilog;
use verilog.vl_types.all;
entity cacheDatapath_sv_unit is
end cacheDatapath_sv_unit;
