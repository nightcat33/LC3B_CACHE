library verilog;
use verilog.vl_types.all;
entity CPU is
end CPU;
