library verilog;
use verilog.vl_types.all;
entity cacheControl_sv_unit is
end cacheControl_sv_unit;
